module filestore

pub struct Disk {
	folder string [required]
}
