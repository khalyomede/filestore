module filestorage

pub struct Disk {
	folder string [required]
}
